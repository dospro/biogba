module biogba